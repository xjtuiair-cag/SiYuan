package swf_pkg;
`include "glb_def.svh"
`include "sy_ovall.svh"
`include "sy_ppl.svh"
`include "sy_cache.svh"
`include "sy_mmu.svh"
endpackage
