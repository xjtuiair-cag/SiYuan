`define VC707
`define PLATFORM_XILINX