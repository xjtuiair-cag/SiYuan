`define GENESYS2
`define PLATFORM_XILINX